*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLY_TEMP_SENS_lpe.spi
#else
.include ../../../work/xsch/RPLY_TEMP_SENS.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}


*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0    dc 0
VDD  VDD  VSS  dc 1.8


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD VSS out RPLY_TEMP_SENS

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(VDD) v(VSS) v(out)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit


#ifdef Debug
dc TEMP -50 100 1
*quit
#else
dc TEMP -50 100 1
write
quit
#endif

.endc

.end
